// Code your design here
// Code your design here
`include "alu.sv"
`include "Control.sv"
`include "dat_mem.sv"
`include "instr_ROM.sv"
//`include "mach_code.txt"
//`include "milestone2_quicktest.sv"
`include "PC.sv"
`include "PC_LUT.sv"
//`include "prog3.sv"
`include "reg_file.sv"
`include "top_level.sv"
